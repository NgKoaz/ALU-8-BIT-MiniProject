module adder_8bit(
    input [7:0] a,
    input [7:0] b,
    input c_in,
    output [8:0] sum,
    output c_out,
);

    // Concate 8 full adder add here
    


endmodule
